package base_pkg;
    typedef logic [31:0] data_32_t;
    typedef logic [15:0] addr_16_t;
    typedef logic [3:0] mask4_t;
endpackage