interface data_transfer;
    
    logic [7:0] mdata;
    logic [7:0] sdata;

endinterface 